library IEEE;
use IEEE.STD_LOGIC_1164.ALL;

entity FF_D16 is
    port (
        clk   : in  std_logic;
        rst_n : in  std_logic;
        d     : in  std_logic_vector(15 downto 0);
        q     : out std_logic_vector(15 downto 0)
    );
end entity;

architecture rtl of FF_D16 is
begin
    process (clk, rst_n)
    begin
        if rst_n = '0' then
            q <= (others => '0');
        elsif rising_edge(clk) then
            q <= d;
        end if;
    end process;
end architecture;